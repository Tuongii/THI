	LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.all;
	USE IEEE.STD_LOGIC_ARITH.ALL;
	USE IEEE.STD_LOGIC_UNSIGNED.ALL;
	
	ENTITY D_FF IS 
		PORT(
			SET,CLR	:	IN	STD_LOGIC;
			CLK		:	IN  STD_LOGIC;
			D 		:   IN STD_LOGIC;
			Q 		:   OUT STD_LOGIC;
			NQ 		:   OUT STD_LOGIC
		);
	END ENTITY;

	ARCHITECTURE BEHAVIORAL OF D_FF IS 
		SIGNAL Q1 : STD_LOGIC;
		BEGIN 
			PROCESS(CLK,SET,CLR,D)
				BEGIN
					IF SET ='0' AND CLR ='1' THEN Q1 <='1';
					ELSIF SET='1' AND CLR ='1' THEN Q1 <='0';
					ELSIF SET ='1' AND CLR ='1' THEN
						IF RISING_EDGE(CLK) THEN
							IF D='1' THEN Q1 <='1';
							ELSIF D ='0' THEN Q1 <='0';
							END IF;
						END IF;
					END IF;
			END PROCESS;
			Q <= Q1;
			NQ <= NOT Q1;

	END BEHAVIORAL;
			